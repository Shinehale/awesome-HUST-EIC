`timescale 1ns / 1ps
module T_4_16(A, EN, Q);
input EN;
input [3:0] A;
output wire [15:0] Q;

reg [15: 0] qregs;

always @(*) begin
    if (EN == 1'b1) begin
        case(A[3:0])
            4'b0000: qregs[15:0] <= 16'b0000000000000001;
            4'b0001: qregs[15:0] <= 16'b0000000000000010;
            4'b0010: qregs[15:0] <= 16'b0000000000000100;
            4'b0011: qregs[15:0] <= 16'b0000000000001000;
            4'b0100: qregs[15:0] <= 16'b0000000000010000;
            4'b0101: qregs[15:0] <= 16'b0000000000100000;
            4'b0110: qregs[15:0] <= 16'b0000000001000000;
            4'b0111: qregs[15:0] <= 16'b0000000010000000;
            4'b1000: qregs[15:0] <= 16'b0000000100000000;
            4'b1001: qregs[15:0] <= 16'b0000001000000000;
            4'b1010: qregs[15:0] <= 16'b0000010000000000;
            4'b1011: qregs[15:0] <= 16'b0000100000000000;
            4'b1100: qregs[15:0] <= 16'b0001000000000000;
            4'b1101: qregs[15:0] <= 16'b0010000000000000;
            4'b1110: qregs[15:0] <= 16'b0100000000000000;
            4'b1111: qregs[15:0] <= 16'b1000000000000000;
	endcase
    end

    else begin
        qregs[15:0] <= 16'b0000000000000000;
    end
end
 
assign Q = qregs;

endmodule
